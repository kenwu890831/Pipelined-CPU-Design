
module Shifter( inputNum, move, Signal , dataOut );

input [31:0]  inputNum ;
input [31:0]  move ;
input [5:0]  Signal  ;
output [31:0] dataOut ;
input reset ;
reg [31:0] zero = 32'b0;
reg [5:0] ctrl = 6'b100000;
reg [31:0] temp =32'b0 ;
parameter SLL = 6'b000000;

wire [31:0] saveOne ;
wire [31:0] saveTwo ;
wire [31:0] saveThree ;
wire [31:0] saveFour ;
wire [31:0] saveFive ;


//16bit 
Shifter_mux2x1  ins_431 ( inputNum[31], inputNum[15], move[4], saveOne[31], Signal );
Shifter_mux2x1  ins_430 ( inputNum[30], inputNum[14], move[4], saveOne[30], Signal );
Shifter_mux2x1  ins_429 ( inputNum[29], inputNum[13], move[4], saveOne[29], Signal );
Shifter_mux2x1  ins_428 ( inputNum[28], inputNum[12], move[4], saveOne[28], Signal );
Shifter_mux2x1  ins_427 ( inputNum[27], inputNum[11], move[4], saveOne[27], Signal );
Shifter_mux2x1  ins_426 ( inputNum[26], inputNum[10], move[4], saveOne[26], Signal );
Shifter_mux2x1  ins_425 ( inputNum[25], inputNum[9], move[4], saveOne[25], Signal );
Shifter_mux2x1  ins_424 ( inputNum[24], inputNum[8], move[4], saveOne[24], Signal );
Shifter_mux2x1  ins_423 ( inputNum[23], inputNum[7], move[4], saveOne[23], Signal );
Shifter_mux2x1  ins_422 ( inputNum[22], inputNum[6], move[4], saveOne[22], Signal );
Shifter_mux2x1  ins_421 ( inputNum[21], inputNum[5], move[4], saveOne[21], Signal );
Shifter_mux2x1  ins_420 ( inputNum[20], inputNum[4], move[4], saveOne[20], Signal );
Shifter_mux2x1  ins_419 ( inputNum[19], inputNum[3], move[4], saveOne[19], Signal );
Shifter_mux2x1  ins_418 ( inputNum[18], inputNum[2], move[4], saveOne[18], Signal );
Shifter_mux2x1  ins_417 ( inputNum[17], inputNum[1], move[4], saveOne[17], Signal );
Shifter_mux2x1  ins_416 ( inputNum[16], inputNum[0], move[4], saveOne[16], Signal );
Shifter_mux2x1  ins_415 ( inputNum[15],1'b0, move[4], saveOne[15], Signal );
Shifter_mux2x1  ins_414 ( inputNum[14],1'b0, move[4], saveOne[14], Signal );
Shifter_mux2x1  ins_413 ( inputNum[13],1'b0, move[4], saveOne[13], Signal );
Shifter_mux2x1  ins_412 ( inputNum[12],1'b0, move[4], saveOne[12], Signal );
Shifter_mux2x1  ins_411 ( inputNum[11],1'b0, move[4], saveOne[11], Signal );
Shifter_mux2x1  ins_410 ( inputNum[10],1'b0, move[4], saveOne[10], Signal );
Shifter_mux2x1  ins_409 ( inputNum[9],1'b0, move[4], saveOne[9], Signal );
Shifter_mux2x1  ins_408 ( inputNum[8],1'b0, move[4], saveOne[8], Signal );
Shifter_mux2x1  ins_407 ( inputNum[7],1'b0, move[4], saveOne[7], Signal );
Shifter_mux2x1  ins_406 ( inputNum[6],1'b0, move[4], saveOne[6], Signal );
Shifter_mux2x1  ins_405 ( inputNum[5],1'b0, move[4], saveOne[5], Signal );
Shifter_mux2x1  ins_404 ( inputNum[4],1'b0, move[4], saveOne[4], Signal );
Shifter_mux2x1  ins_403 ( inputNum[3],1'b0, move[4], saveOne[3], Signal );
Shifter_mux2x1  ins_402 ( inputNum[2],1'b0, move[4], saveOne[2], Signal );
Shifter_mux2x1  ins_401 ( inputNum[1],1'b0, move[4], saveOne[1], Signal );
Shifter_mux2x1  ins_400 ( inputNum[0],1'b0, move[4], saveOne[0], Signal );

//8bit
Shifter_mux2x1  ins_331 ( saveOne[31], saveOne[23], move[3], saveTwo[31], Signal );
Shifter_mux2x1  ins_330 ( saveOne[30], saveOne[22], move[3], saveTwo[30], Signal );
Shifter_mux2x1  ins_329 ( saveOne[29], saveOne[21], move[3], saveTwo[29], Signal );
Shifter_mux2x1  ins_328 ( saveOne[28], saveOne[20], move[3], saveTwo[28], Signal );
Shifter_mux2x1  ins_327 ( saveOne[27], saveOne[19], move[3], saveTwo[27], Signal );
Shifter_mux2x1  ins_326 ( saveOne[26], saveOne[18], move[3], saveTwo[26], Signal );
Shifter_mux2x1  ins_325 ( saveOne[25], saveOne[17], move[3], saveTwo[25], Signal );
Shifter_mux2x1  ins_324 ( saveOne[24], saveOne[16], move[3], saveTwo[24], Signal );
Shifter_mux2x1  ins_323 ( saveOne[23], saveOne[15], move[3], saveTwo[23], Signal );
Shifter_mux2x1  ins_322 ( saveOne[22], saveOne[14], move[3], saveTwo[22], Signal );
Shifter_mux2x1  ins_321 ( saveOne[21], saveOne[13], move[3], saveTwo[21], Signal );
Shifter_mux2x1  ins_320 ( saveOne[20], saveOne[12], move[3], saveTwo[20], Signal );
Shifter_mux2x1  ins_319 ( saveOne[19], saveOne[11], move[3], saveTwo[19], Signal );
Shifter_mux2x1  ins_318 ( saveOne[18], saveOne[10], move[3], saveTwo[18], Signal );
Shifter_mux2x1  ins_317 ( saveOne[17], saveOne[9], move[3], saveTwo[17], Signal );
Shifter_mux2x1  ins_316 ( saveOne[16], saveOne[8], move[3], saveTwo[16], Signal );
Shifter_mux2x1  ins_315 ( saveOne[15], saveOne[7], move[3], saveTwo[15], Signal );
Shifter_mux2x1  ins_314 ( saveOne[14], saveOne[6], move[3], saveTwo[14], Signal );
Shifter_mux2x1  ins_313 ( saveOne[13], saveOne[5], move[3], saveTwo[13], Signal );
Shifter_mux2x1  ins_312 ( saveOne[12], saveOne[4], move[3], saveTwo[12], Signal );
Shifter_mux2x1  ins_311 ( saveOne[11], saveOne[3], move[3], saveTwo[11], Signal );
Shifter_mux2x1  ins_310 ( saveOne[10], saveOne[2], move[3], saveTwo[10], Signal );
Shifter_mux2x1  ins_309 ( saveOne[9], saveOne[1], move[3], saveTwo[9], Signal );
Shifter_mux2x1  ins_308 ( saveOne[8], saveOne[0], move[3], saveTwo[8], Signal );
Shifter_mux2x1  ins_307 ( saveOne[7],1'b0, move[3], saveTwo[7], Signal );
Shifter_mux2x1  ins_306 ( saveOne[6],1'b0, move[3], saveTwo[6], Signal );
Shifter_mux2x1  ins_305 ( saveOne[5],1'b0, move[3], saveTwo[5], Signal );
Shifter_mux2x1  ins_304 ( saveOne[4],1'b0, move[3], saveTwo[4], Signal );
Shifter_mux2x1  ins_303 ( saveOne[3],1'b0, move[3], saveTwo[3], Signal );
Shifter_mux2x1  ins_302 ( saveOne[2],1'b0, move[3], saveTwo[2], Signal );
Shifter_mux2x1  ins_301 ( saveOne[1],1'b0, move[3], saveTwo[1], Signal );
Shifter_mux2x1  ins_300 ( saveOne[0],1'b0, move[3], saveTwo[0], Signal );

//4bit 
Shifter_mux2x1  ins_231 ( saveTwo[31], saveTwo[27], move[2], saveThree[31], Signal );
Shifter_mux2x1  ins_230 ( saveTwo[30], saveTwo[26], move[2], saveThree[30], Signal );
Shifter_mux2x1  ins_229 ( saveTwo[29], saveTwo[25], move[2], saveThree[29], Signal );
Shifter_mux2x1  ins_228 ( saveTwo[28], saveTwo[24], move[2], saveThree[28], Signal );
Shifter_mux2x1  ins_227 ( saveTwo[27], saveTwo[23], move[2], saveThree[27], Signal );
Shifter_mux2x1  ins_226 ( saveTwo[26], saveTwo[22], move[2], saveThree[26], Signal );
Shifter_mux2x1  ins_225 ( saveTwo[25], saveTwo[21], move[2], saveThree[25], Signal );
Shifter_mux2x1  ins_224 ( saveTwo[24], saveTwo[20], move[2], saveThree[24], Signal );
Shifter_mux2x1  ins_223 ( saveTwo[23], saveTwo[19], move[2], saveThree[23], Signal );
Shifter_mux2x1  ins_222 ( saveTwo[22], saveTwo[18], move[2], saveThree[22], Signal );
Shifter_mux2x1  ins_221 ( saveTwo[21], saveTwo[17], move[2], saveThree[21], Signal );
Shifter_mux2x1  ins_220 ( saveTwo[20], saveTwo[16], move[2], saveThree[20], Signal );
Shifter_mux2x1  ins_219 ( saveTwo[19], saveTwo[15], move[2], saveThree[19], Signal );
Shifter_mux2x1  ins_218 ( saveTwo[18], saveTwo[14], move[2], saveThree[18], Signal );
Shifter_mux2x1  ins_217 ( saveTwo[17], saveTwo[13], move[2], saveThree[17], Signal );
Shifter_mux2x1  ins_216 ( saveTwo[16], saveTwo[12], move[2], saveThree[16], Signal );
Shifter_mux2x1  ins_215 ( saveTwo[15], saveTwo[11], move[2], saveThree[15], Signal );
Shifter_mux2x1  ins_214 ( saveTwo[14], saveTwo[10], move[2], saveThree[14], Signal );
Shifter_mux2x1  ins_213 ( saveTwo[13], saveTwo[9], move[2], saveThree[13], Signal );
Shifter_mux2x1  ins_212 ( saveTwo[12], saveTwo[8], move[2], saveThree[12], Signal );
Shifter_mux2x1  ins_211 ( saveTwo[11], saveTwo[7], move[2], saveThree[11], Signal );
Shifter_mux2x1  ins_210 ( saveTwo[10], saveTwo[6], move[2], saveThree[10], Signal );
Shifter_mux2x1  ins_209 ( saveTwo[9], saveTwo[5], move[2], saveThree[9], Signal );
Shifter_mux2x1  ins_208 ( saveTwo[8], saveTwo[4], move[2], saveThree[8], Signal );
Shifter_mux2x1  ins_207 ( saveTwo[7], saveTwo[3], move[2], saveThree[7], Signal );
Shifter_mux2x1  ins_206 ( saveTwo[6], saveTwo[2], move[2], saveThree[6], Signal );
Shifter_mux2x1  ins_205 ( saveTwo[5], saveTwo[1], move[2], saveThree[5], Signal );
Shifter_mux2x1  ins_204 ( saveTwo[4], saveTwo[0], move[2], saveThree[4], Signal );
Shifter_mux2x1  ins_203 ( saveTwo[3],1'b0, move[2], saveThree[3], Signal );
Shifter_mux2x1  ins_202 ( saveTwo[2],1'b0, move[2], saveThree[2], Signal );
Shifter_mux2x1  ins_201 ( saveTwo[1],1'b0, move[2], saveThree[1], Signal );
Shifter_mux2x1  ins_200 ( saveTwo[0],1'b0, move[2], saveThree[0], Signal );

// 2 bit
Shifter_mux2x1  ins_131 ( saveThree[31], saveThree[29], move[1], saveFour[31], Signal );
Shifter_mux2x1  ins_130 ( saveThree[30], saveThree[28], move[1], saveFour[30], Signal );
Shifter_mux2x1  ins_129 ( saveThree[29], saveThree[27], move[1], saveFour[29], Signal );
Shifter_mux2x1  ins_128 ( saveThree[28], saveThree[26], move[1], saveFour[28], Signal );
Shifter_mux2x1  ins_127 ( saveThree[27], saveThree[25], move[1], saveFour[27], Signal );
Shifter_mux2x1  ins_126 ( saveThree[26], saveThree[24], move[1], saveFour[26], Signal );
Shifter_mux2x1  ins_125 ( saveThree[25], saveThree[23], move[1], saveFour[25], Signal );
Shifter_mux2x1  ins_124 ( saveThree[24], saveThree[22], move[1], saveFour[24], Signal );
Shifter_mux2x1  ins_123 ( saveThree[23], saveThree[21], move[1], saveFour[23], Signal );
Shifter_mux2x1  ins_122 ( saveThree[22], saveThree[20], move[1], saveFour[22], Signal );
Shifter_mux2x1  ins_121 ( saveThree[21], saveThree[19], move[1], saveFour[21], Signal );
Shifter_mux2x1  ins_120 ( saveThree[20], saveThree[18], move[1], saveFour[20], Signal );
Shifter_mux2x1  ins_119 ( saveThree[19], saveThree[17], move[1], saveFour[19], Signal );
Shifter_mux2x1  ins_118 ( saveThree[18], saveThree[16], move[1], saveFour[18], Signal );
Shifter_mux2x1  ins_117 ( saveThree[17], saveThree[15], move[1], saveFour[17], Signal );
Shifter_mux2x1  ins_116 ( saveThree[16], saveThree[14], move[1], saveFour[16], Signal );
Shifter_mux2x1  ins_115 ( saveThree[15], saveThree[13], move[1], saveFour[15], Signal );
Shifter_mux2x1  ins_114 ( saveThree[14], saveThree[12], move[1], saveFour[14], Signal );
Shifter_mux2x1  ins_113 ( saveThree[13], saveThree[11], move[1], saveFour[13], Signal );
Shifter_mux2x1  ins_112 ( saveThree[12], saveThree[10], move[1], saveFour[12], Signal );
Shifter_mux2x1  ins_111 ( saveThree[11], saveThree[9], move[1], saveFour[11], Signal );
Shifter_mux2x1  ins_110 ( saveThree[10], saveThree[8], move[1], saveFour[10], Signal );
Shifter_mux2x1  ins_109 ( saveThree[9], saveThree[7], move[1], saveFour[9], Signal );
Shifter_mux2x1  ins_108 ( saveThree[8], saveThree[6], move[1], saveFour[8], Signal );
Shifter_mux2x1  ins_107 ( saveThree[7], saveThree[5], move[1], saveFour[7], Signal );
Shifter_mux2x1  ins_106 ( saveThree[6], saveThree[4], move[1], saveFour[6], Signal );
Shifter_mux2x1  ins_105 ( saveThree[5], saveThree[3], move[1], saveFour[5], Signal );
Shifter_mux2x1  ins_104 ( saveThree[4], saveThree[2], move[1], saveFour[4], Signal );
Shifter_mux2x1  ins_103 ( saveThree[3], saveThree[1], move[1], saveFour[3], Signal );
Shifter_mux2x1  ins_102 ( saveThree[2], saveThree[0], move[1], saveFour[2], Signal );
Shifter_mux2x1  ins_101 ( saveThree[1],1'b0, move[1], saveFour[1], Signal );
Shifter_mux2x1  ins_100 ( saveThree[0],1'b0, move[1], saveFour[0], Signal );

// bit1
Shifter_mux2x1  ins_031 ( saveFour[31], saveFour[30], move[0], saveFive[31], Signal );
Shifter_mux2x1  ins_030 ( saveFour[30], saveFour[29], move[0], saveFive[30], Signal );
Shifter_mux2x1  ins_029 ( saveFour[29], saveFour[28], move[0], saveFive[29], Signal );
Shifter_mux2x1  ins_028 ( saveFour[28], saveFour[27], move[0], saveFive[28], Signal );
Shifter_mux2x1  ins_027 ( saveFour[27], saveFour[26], move[0], saveFive[27], Signal );
Shifter_mux2x1  ins_026 ( saveFour[26], saveFour[25], move[0], saveFive[26], Signal );
Shifter_mux2x1  ins_025 ( saveFour[25], saveFour[24], move[0], saveFive[25], Signal );
Shifter_mux2x1  ins_024 ( saveFour[24], saveFour[23], move[0], saveFive[24], Signal );
Shifter_mux2x1  ins_023 ( saveFour[23], saveFour[22], move[0], saveFive[23], Signal );
Shifter_mux2x1  ins_022 ( saveFour[22], saveFour[21], move[0], saveFive[22], Signal );
Shifter_mux2x1  ins_021 ( saveFour[21], saveFour[20], move[0], saveFive[21], Signal );
Shifter_mux2x1  ins_020 ( saveFour[20], saveFour[19], move[0], saveFive[20], Signal );
Shifter_mux2x1  ins_019 ( saveFour[19], saveFour[18], move[0], saveFive[19], Signal );
Shifter_mux2x1  ins_018 ( saveFour[18], saveFour[17], move[0], saveFive[18], Signal );
Shifter_mux2x1  ins_017 ( saveFour[17], saveFour[16], move[0], saveFive[17], Signal );
Shifter_mux2x1  ins_016 ( saveFour[16], saveFour[15], move[0], saveFive[16], Signal );
Shifter_mux2x1  ins_015 ( saveFour[15], saveFour[14], move[0], saveFive[15], Signal );
Shifter_mux2x1  ins_014 ( saveFour[14], saveFour[13], move[0], saveFive[14], Signal );
Shifter_mux2x1  ins_013 ( saveFour[13], saveFour[12], move[0], saveFive[13], Signal );
Shifter_mux2x1  ins_012 ( saveFour[12], saveFour[11], move[0], saveFive[12], Signal );
Shifter_mux2x1  ins_011 ( saveFour[11], saveFour[10], move[0], saveFive[11], Signal );
Shifter_mux2x1  ins_010 ( saveFour[10], saveFour[9], move[0], saveFive[10], Signal );
Shifter_mux2x1  ins_009 ( saveFour[9], saveFour[8], move[0], saveFive[9], Signal );
Shifter_mux2x1  ins_008 ( saveFour[8], saveFour[7], move[0], saveFive[8], Signal );
Shifter_mux2x1  ins_007 ( saveFour[7], saveFour[6], move[0], saveFive[7], Signal );
Shifter_mux2x1  ins_006 ( saveFour[6], saveFour[5], move[0], saveFive[6], Signal );
Shifter_mux2x1  ins_005 ( saveFour[5], saveFour[4], move[0], saveFive[5], Signal );
Shifter_mux2x1  ins_004 ( saveFour[4], saveFour[3], move[0], saveFive[4], Signal );
Shifter_mux2x1  ins_003 ( saveFour[3], saveFour[2], move[0], saveFive[3], Signal );
Shifter_mux2x1  ins_002 ( saveFour[2], saveFour[1], move[0], saveFive[2], Signal );
Shifter_mux2x1  ins_001 ( saveFour[1], saveFour[0], move[0], saveFive[1], Signal );
Shifter_mux2x1  ins_000 ( saveFour[0],1'b0, move[0], saveFive[0], Signal );

assign dataOut = ( move >= ctrl)? zero : saveFive ;

endmodule
